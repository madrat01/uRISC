module top_tb();

logic clk;
logic rst;
logic err;

top uRISC(.*);

endmodule